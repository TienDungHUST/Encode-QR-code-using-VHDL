library verilog;
use verilog.vl_types.all;
entity test_xor_int_vlg_vec_tst is
end test_xor_int_vlg_vec_tst;
