library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
--USE work.data_types.all; 
------------------------------------
package my_package is
TYPE my_integer IS RANGE 0 to 255;
	function Convert_to_anpha(inte : in my_integer) return my_integer;
	function Convert_to_integer(inte : in my_integer) return my_integer;

end package my_package;
------------------------------------
package body my_package is
	function Convert_to_anpha(inte : in my_integer) return my_integer;
	function Convert_to_integer(anpha : in my_integer) return my_integer;
-- Function convert integer totemp2 
FUNCTION Convert_to_anpha(inte : in my_integer) return my_integer IS
	variable temp1 : INTEGER;
BEGIN
	CASE inte IS
		WHEN 1 => temp1 := 0 ;
		WHEN 2 => temp1 := 1 ;
		WHEN 3 => temp1 := 25 ;
		WHEN 4 => temp1 := 2 ;
		WHEN 5 => temp1 := 50 ;
		WHEN 6 => temp1 := 26 ;
		WHEN 7 => temp1 := 198 ;
		WHEN 8 => temp1 := 3 ;
		WHEN 9 => temp1 := 223 ;
		WHEN 10 => temp1 := 51 ;
		WHEN 11 => temp1 := 238 ;
		WHEN 12 => temp1 := 27 ;
		WHEN 13 => temp1 := 104 ;
		WHEN 14 => temp1 := 199 ;
		WHEN 15 => temp1 := 75 ;
		WHEN 16 => temp1 := 4 ;
		WHEN 17 => temp1 := 100 ;
		WHEN 18 => temp1 := 224 ;
		WHEN 19 => temp1 := 14 ;
		WHEN 20 => temp1 := 52 ;
		WHEN 21 => temp1 := 141 ;
		WHEN 22 => temp1 := 239 ;
		WHEN 23 => temp1 := 129 ;
		WHEN 24 => temp1 := 28 ;
		WHEN 25 => temp1 := 193 ;
		WHEN 26 => temp1 := 105 ;
		WHEN 27 => temp1 := 248 ;
		WHEN 28 => temp1 := 200 ;
		WHEN 29 => temp1 := 8 ;
		WHEN 30 => temp1 := 76 ;
		WHEN 31 => temp1 := 113 ;
		WHEN 32 => temp1 := 5 ;
		WHEN 33 => temp1 := 138 ;
		WHEN 34 => temp1 := 101 ;
		WHEN 35 => temp1 := 47 ;
		WHEN 36 => temp1 := 225 ;
		WHEN 37 => temp1 := 36 ;
		WHEN 38 => temp1 := 15 ;
		WHEN 39 => temp1 := 33 ;
		WHEN 40 => temp1 := 53 ;
		WHEN 41 => temp1 := 147 ;
		WHEN 42 => temp1 := 142 ;
		WHEN 43 => temp1 := 218 ;
		WHEN 44 => temp1 := 240 ;
		WHEN 45 => temp1 := 18 ;
		WHEN 46 => temp1 := 130 ;
		WHEN 47 => temp1 := 69 ;
		WHEN 48 => temp1 := 29 ;
		WHEN 49 => temp1 := 181 ;
		WHEN 50 => temp1 := 194 ;
		WHEN 51 => temp1 := 125 ;
		WHEN 52 => temp1 := 106 ;
		WHEN 53 => temp1 := 39 ;
		WHEN 54 => temp1 := 249 ;
		WHEN 55 => temp1 := 185 ;
		WHEN 56 => temp1 := 201 ;
		WHEN 57 => temp1 := 154 ;
		WHEN 58 => temp1 := 9 ;
		WHEN 59 => temp1 := 120 ;
		WHEN 60 => temp1 := 77 ;
		WHEN 61 => temp1 := 228 ;
		WHEN 62 => temp1 := 114 ;
		WHEN 63 => temp1 := 166 ;
		WHEN 64 => temp1 := 6 ;
		WHEN 65 => temp1 := 191 ;
		WHEN 66 => temp1 := 139 ;
		WHEN 67 => temp1 := 98 ;
		WHEN 68 => temp1 := 102 ;
		WHEN 69 => temp1 := 221 ;
		WHEN 70 => temp1 := 48 ;
		WHEN 71 => temp1 := 253 ;
		WHEN 72 => temp1 := 226 ;
		WHEN 73 => temp1 := 152 ;
		WHEN 74 => temp1 := 37 ;
		WHEN 75 => temp1 := 179 ;
		WHEN 76 => temp1 := 16 ;
		WHEN 77 => temp1 := 145 ;
		WHEN 78 => temp1 := 34 ;
		WHEN 79 => temp1 := 136 ;
		WHEN 80 => temp1 := 54 ;
		WHEN 81 => temp1 := 208 ;
		WHEN 82 => temp1 := 148 ;
		WHEN 83 => temp1 := 206 ;
		WHEN 84 => temp1 := 143 ;
		WHEN 85 => temp1 := 150 ;
		WHEN 86 => temp1 := 219 ;
		WHEN 87 => temp1 := 189 ;
		WHEN 88 => temp1 := 241 ;
		WHEN 89 => temp1 := 210 ;
		WHEN 90 => temp1 := 19 ;
		WHEN 91 => temp1 := 92 ;
		WHEN 92 => temp1 := 131 ;
		WHEN 93 => temp1 := 56 ;
		WHEN 94 => temp1 := 70 ;
		WHEN 95 => temp1 := 64 ;
		WHEN 96 => temp1 := 30 ;
		WHEN 97 => temp1 := 66 ;
		WHEN 98 => temp1 := 182 ;
		WHEN 99 => temp1 := 163 ;
		WHEN 100 => temp1 := 195 ;
		WHEN 101 => temp1 := 72 ;
		WHEN 102 => temp1 := 126;
		WHEN 103 => temp1 := 110 ;
		WHEN 104 => temp1 := 107 ;
		WHEN 105 => temp1 := 58 ;
		WHEN 106 => temp1 := 40 ;
		WHEN 107 => temp1 := 84 ;
		WHEN 108 => temp1 := 250 ;
		WHEN 109 => temp1 := 133 ;
		WHEN 110 => temp1 := 186 ;
		WHEN 111 => temp1 := 61 ;
		WHEN 112 => temp1 := 202 ;
		WHEN 113 => temp1 := 94 ;
		WHEN 114 => temp1 := 155 ;
		WHEN 115 => temp1 := 159 ;
		WHEN 116 => temp1 := 10 ;
		WHEN 117 => temp1 := 21 ;
		WHEN 118 => temp1 := 121 ;
		WHEN 119 => temp1 := 43 ;
		WHEN 120 => temp1 := 78 ;
		WHEN 121 => temp1 := 212 ;
		WHEN 122 => temp1 := 229 ;
		WHEN 123 => temp1 := 172 ;
		WHEN 124 => temp1 := 115 ;
		WHEN 125 => temp1 := 243 ;
		WHEN 126 => temp1 := 167 ;
		WHEN 127 => temp1 := 87 ;
		WHEN 128 => temp1 := 7 ;
		WHEN 129 => temp1 := 112 ;
		WHEN 130 => temp1 := 192 ;
		WHEN 131 => temp1 := 247 ;
		WHEN 132 => temp1 := 140 ;
		WHEN 133 => temp1 := 128 ;
		WHEN 134 => temp1 := 99 ;
		WHEN 135 => temp1 := 13 ;
		WHEN 136 => temp1 := 103 ;
		WHEN 137 => temp1 := 74 ;
		WHEN 138 => temp1 := 222 ;
		WHEN 139 => temp1 := 237 ;
		WHEN 140 => temp1 := 49 ;
		WHEN 141 => temp1 := 197 ;
		WHEN 142 => temp1 := 254 ;
		WHEN 143 => temp1 := 24 ;
		WHEN 144 => temp1 := 227 ;
		WHEN 145 => temp1 := 165 ;
		WHEN 146 => temp1 := 153 ;
		WHEN 147 => temp1 := 119 ;
		WHEN 148 => temp1 := 38 ;
		WHEN 149 => temp1 := 184 ;
		WHEN 150 => temp1 := 180 ;
		WHEN 151 => temp1 := 124 ;
		WHEN 152 => temp1 := 17 ;
		WHEN 153 => temp1 := 68 ;
		WHEN 154 => temp1 := 146 ;
		WHEN 155 => temp1 := 217 ;
		WHEN 156 => temp1 := 35 ;
		WHEN 157 => temp1 := 32 ;
		WHEN 158 => temp1 := 137 ;
		WHEN 159 => temp1 := 46 ;
		WHEN 160 => temp1 := 55 ;
		WHEN 161 => temp1 := 63 ;
		WHEN 162 => temp1 := 209 ;
		WHEN 163 => temp1 := 91 ;
		WHEN 164 => temp1 := 149 ;
		WHEN 165 => temp1 := 188 ;
		WHEN 166 => temp1 := 207 ;
		WHEN 167 => temp1 := 205 ;
		WHEN 168 => temp1 := 144 ;
		WHEN 169 => temp1 := 135 ;
		WHEN 170 => temp1 := 151 ;
		WHEN 171 => temp1 := 178 ;
		WHEN 172 => temp1 := 220 ;
		WHEN 173 => temp1 := 252 ;
		WHEN 174 => temp1 := 190 ;
		WHEN 175 => temp1 := 97 ;
		WHEN 176 => temp1 := 242;
		WHEN 177 => temp1 := 86 ;
		WHEN 178 => temp1 := 211 ;
		WHEN 179 => temp1 := 171 ;
		WHEN 180 => temp1 := 20 ;
		WHEN 181 => temp1 := 42 ;
		WHEN 182 => temp1 := 93 ;
		WHEN 183 => temp1 := 158 ;
		WHEN 184 => temp1 := 132 ;
		WHEN 185 => temp1 := 60 ;
		WHEN 186 => temp1 := 57 ;
		WHEN 187 => temp1 := 83 ;
		WHEN 188 => temp1 := 71 ;
		WHEN 189 => temp1 := 109 ;
		WHEN 190 => temp1 := 65 ;
		WHEN 191 => temp1 := 162;
		WHEN 192 => temp1 := 31 ;
		WHEN 193 => temp1 := 45 ;
		WHEN 194 => temp1 := 67 ;
		WHEN 195 => temp1 := 216 ;
		WHEN 196 => temp1 := 183 ;
		WHEN 197 => temp1 := 123 ;
		WHEN 198 => temp1 := 164 ;
		WHEN 199 => temp1 := 118;
		WHEN 200 => temp1 := 196 ;
		WHEN 201 => temp1 := 23 ;
		WHEN 202 => temp1 := 73 ;
		WHEN 203 => temp1 := 236 ;
		WHEN 204 => temp1 := 127 ;
		WHEN 205 => temp1 := 12 ;
		WHEN 206 => temp1 := 111 ;
		WHEN 207 => temp1 := 246 ;
		WHEN 208 => temp1 := 108 ;
		WHEN 209 => temp1 := 161 ;
		WHEN 210 => temp1 := 59 ;
		WHEN 211 => temp1 := 82 ;
		WHEN 212 => temp1 := 41 ;
		WHEN 213 => temp1 := 157 ;
		WHEN 214 => temp1 := 85 ;
		WHEN 215 => temp1 := 170 ;
		WHEN 216 => temp1 := 251 ;
		WHEN 217 => temp1 := 96 ;
		WHEN 218 => temp1 := 134 ;
		WHEN 219 => temp1 := 177 ;
		WHEN 220 => temp1 := 187 ;
		WHEN 221 => temp1 := 204 ;
		WHEN 222 => temp1 := 62 ;
		WHEN 223 => temp1 := 90 ;
		WHEN 224 => temp1 := 203 ;
		WHEN 225 => temp1 := 89 ;
		WHEN 226 => temp1 := 95 ;
		WHEN 227 => temp1 := 176 ;
		WHEN 228 => temp1 := 156 ;
		WHEN 229 => temp1 := 169 ;
		WHEN 230 => temp1 := 160 ;
		WHEN 231 => temp1 := 81 ;
		WHEN 232 => temp1 := 11 ;
		WHEN 233 => temp1 := 245 ;
		WHEN 234 => temp1 := 22 ;
		WHEN 235 => temp1 := 235 ;
		WHEN 236 => temp1 := 122 ;
		WHEN 237 => temp1 := 117 ;
		WHEN 238 => temp1 := 44 ;
		WHEN 239 => temp1 := 215 ;
		WHEN 240 => temp1 := 79 ;
		WHEN 241 => temp1 := 174 ;
		WHEN 242 => temp1 := 213 ;
		WHEN 243 => temp1 := 233 ;
		WHEN 244 => temp1 := 230 ;
		WHEN 245 => temp1 := 231 ;
		WHEN 246 => temp1 := 173 ;
		WHEN 247 => temp1 := 232 ;
		WHEN 248 => temp1 := 116 ;
		WHEN 249 => temp1 := 214 ;
		WHEN 250 => temp1 := 244 ;
		WHEN 251 => temp1 := 234 ;
		WHEN 252 => temp1 := 168 ;
		WHEN 253 => temp1 := 80 ;
		WHEN 254 => temp1 := 88 ;
		WHEN 255 => temp1 := 175 ;
			
		return temp1;
		
		END CASE;
		
END FUNCTION Convert_to_anpha;

--Function convert anphato integer
FUNCTION Convert_to_integer(anpha : in my_integer) return my_integer IS
	variable temp2 : INTEGER RANGE 0 TO 255;
BEGIN
	CASE anpha IS
		WHEN 0 => temp2 := 1 ;
		WHEN 1 => temp2 := 2 ;
		WHEN 2 => temp2 := 4 ;
		WHEN 3 => temp2 := 8 ;
		WHEN 4 => temp2 := 16 ;
		WHEN 5 => temp2 := 32 ;
		WHEN 6 => temp2 := 64 ;
		WHEN 7 => temp2 := 128 ;
		WHEN 8 => temp2 := 29 ;
		WHEN 9 => temp2 := 58 ;
		WHEN 10 => temp2 := 116 ;
		WHEN 11 => temp2 := 232 ;
		WHEN 12 => temp2 := 205 ;
		WHEN 13 => temp2 := 135 ;
		WHEN 14 => temp2 := 19 ;
		WHEN 15 => temp2 := 38 ;
		WHEN 16 => temp2 := 76 ;
		WHEN 17 => temp2 := 152 ;
		WHEN 18 => temp2 := 45 ;
		WHEN 19 => temp2 := 90 ;
		WHEN 20 => temp2 := 180 ;
		WHEN 21 => temp2 := 117 ;
		WHEN 22 => temp2 := 234 ;
		WHEN 23 => temp2 := 201 ;
		WHEN 24 => temp2 := 143 ;
		WHEN 25 => temp2 := 3 ;
		WHEN 26 => temp2 := 6 ;
		WHEN 27 => temp2 := 12 ;
		WHEN 28 => temp2 := 24 ;
		WHEN 29 => temp2 := 48 ;
		WHEN 30 => temp2 := 96 ;
		WHEN 31 => temp2 := 192 ;
		WHEN 32 => temp2 := 157 ;
		WHEN 33 => temp2 := 39 ;
		WHEN 34 => temp2 := 78 ;
		WHEN 35 => temp2 := 156 ;
		WHEN 36 => temp2 := 37 ;
		WHEN 37 => temp2 := 74 ;
		WHEN 38 => temp2 := 148 ;
		WHEN 39 => temp2 := 53 ;
		WHEN 40 => temp2 := 106 ;
		WHEN 41 => temp2 := 212 ;
		WHEN 42 => temp2 := 181 ;
		WHEN 43 => temp2 := 119 ;
		WHEN 44 => temp2 := 238 ;
		WHEN 45 => temp2 := 193 ;
		WHEN 46 => temp2 := 159 ;
		WHEN 47 => temp2 := 35 ;
		WHEN 48 => temp2 := 70 ;
		WHEN 49 => temp2 := 140 ;
		WHEN 50 => temp2 := 5 ;
		WHEN 51 => temp2 := 10 ;
		WHEN 52 => temp2 := 20 ;
		WHEN 53 => temp2 := 40 ;
		WHEN 54 => temp2 := 80 ;
		WHEN 55 => temp2 := 160 ;
		WHEN 56 => temp2 := 93 ;
		WHEN 57 => temp2 := 186 ;
		WHEN 58 => temp2 := 105 ;
		WHEN 59 => temp2 := 210 ;
		WHEN 60 => temp2 := 185 ;
		WHEN 61 => temp2 := 111 ;
		WHEN 62 => temp2 := 222 ;
		WHEN 63 => temp2 := 161 ;
		WHEN 64 => temp2 := 95 ;
		WHEN 65 => temp2 := 190 ;
		WHEN 66 => temp2 := 97 ;
		WHEN 67 => temp2 := 194 ;
		WHEN 68 => temp2 := 153 ;
		WHEN 69 => temp2 := 47 ;
		WHEN 70 => temp2 := 94 ;
		WHEN 71 => temp2 := 188 ;
		WHEN 72 => temp2 := 101 ;
		WHEN 73 => temp2 := 202 ;
		WHEN 74 => temp2 := 137 ;
		WHEN 75 => temp2 := 15 ;
		WHEN 76 => temp2 := 30 ;
		WHEN 77 => temp2 := 60 ;
		WHEN 78 => temp2 := 120 ;
		WHEN 79 => temp2 := 240 ;
		WHEN 80 => temp2 := 253 ;
		WHEN 81 => temp2 := 231 ;
		WHEN 82 => temp2 := 211 ;
		WHEN 83 => temp2 := 187 ;
		WHEN 84 => temp2 := 107 ;
		WHEN 85 => temp2 := 214 ;
		WHEN 86 => temp2 := 177 ;
		WHEN 87 => temp2 := 127 ;
		WHEN 88 => temp2 := 254 ;
		WHEN 89 => temp2 := 225 ;
		WHEN 90 => temp2 := 223 ;
		WHEN 91 => temp2 := 163 ;
		WHEN 92 => temp2 := 91 ;
		WHEN 93 => temp2 := 182 ;
		WHEN 94 => temp2 := 113 ;
		WHEN 95 => temp2 := 226 ;
		WHEN 96 => temp2 := 217 ;
		WHEN 97 => temp2 := 175 ;
		WHEN 98 => temp2 := 67 ;
		WHEN 99 => temp2 := 134 ;
		WHEN 100 => temp2 := 17 ;
		WHEN 101 => temp2 := 34 ;
		WHEN 102 => temp2 := 68 ;
		WHEN 103 => temp2 := 136 ;
		WHEN 104 => temp2 := 13 ;
		WHEN 105 => temp2 := 26 ;
		WHEN 106 => temp2 := 52 ;
		WHEN 107 => temp2 := 104 ;
		WHEN 108 => temp2 := 208 ;
		WHEN 109 => temp2 := 189 ;
		WHEN 110 => temp2 := 103 ;
		WHEN 111 => temp2 := 206 ;
		WHEN 112 => temp2 := 129 ;
		WHEN 113 => temp2 := 31 ;
		WHEN 114 => temp2 := 62 ;
		WHEN 115 => temp2 := 124 ;
		WHEN 116 => temp2 := 248 ;
		WHEN 117 => temp2 := 237 ;
		WHEN 118 => temp2 := 199 ;
		WHEN 119 => temp2 := 147 ;
		WHEN 120 => temp2 := 59 ;
		WHEN 121 => temp2 := 118 ;
		WHEN 122 => temp2 := 236 ;
		WHEN 123 => temp2 := 197 ;
		WHEN 124 => temp2 := 151 ;
		WHEN 125 => temp2 := 51 ;
		WHEN 126 => temp2 := 102 ;
		WHEN 127 => temp2 := 204 ;
		WHEN 128 => temp2 := 133 ;
		WHEN 129 => temp2 := 23 ;
		WHEN 130 => temp2 := 46 ;
		WHEN 131 => temp2 := 92 ;
		WHEN 132 => temp2 := 184 ;
		WHEN 133 => temp2 := 109 ;
		WHEN 134 => temp2 := 218 ;
		WHEN 135 => temp2 := 169 ;
		WHEN 136 => temp2 := 79 ;
		WHEN 137 => temp2 := 158 ;
		WHEN 138 => temp2 := 33 ;
		WHEN 139 => temp2 := 66 ;
		WHEN 140 => temp2 := 132 ;
		WHEN 141 => temp2 := 21 ;
		WHEN 142 => temp2 := 42 ;
		WHEN 143 => temp2 := 84 ;
		WHEN 144 => temp2 := 168 ;
		WHEN 145 => temp2 := 77 ;
		WHEN 146 => temp2 := 154 ;
		WHEN 147 => temp2 := 41 ;
		WHEN 148 => temp2 := 82 ;
		WHEN 149 => temp2 := 164 ;
		WHEN 150 => temp2 := 85 ;
		WHEN 151 => temp2 := 170 ;
		WHEN 152 => temp2 := 73 ;
		WHEN 153 => temp2 := 146 ;
		WHEN 154 => temp2 := 57 ;
		WHEN 155 => temp2 := 114 ;
		WHEN 156 => temp2 := 228 ;
		WHEN 157 => temp2 := 213 ;
		WHEN 158 => temp2 := 183 ;
		WHEN 159 => temp2 := 115 ;
		WHEN 160 => temp2 := 230 ;
		WHEN 161 => temp2 := 209 ;
		WHEN 162 => temp2 := 191 ;
		WHEN 163 => temp2 := 99 ;
		WHEN 164 => temp2 := 198 ;
		WHEN 165 => temp2 := 145 ;
		WHEN 166 => temp2 := 63 ;
		WHEN 167 => temp2 := 126 ;
		WHEN 168 => temp2 := 252 ;
		WHEN 169 => temp2 := 229 ;
		WHEN 170 => temp2 := 215 ;
		WHEN 171 => temp2 := 179 ;
		WHEN 172 => temp2 := 123 ;
		WHEN 173 => temp2 := 246 ;
		WHEN 174 => temp2 := 241 ;
		WHEN 175 => temp2 := 255 ;
		WHEN 176 => temp2 := 227 ;
		WHEN 177 => temp2 := 219 ;
		WHEN 178 => temp2 := 171 ;
		WHEN 179 => temp2 := 75 ;
		WHEN 180 => temp2 := 150 ;
		WHEN 181 => temp2 := 49 ;
		WHEN 182 => temp2 := 98 ;
		WHEN 183 => temp2 := 196 ;
		WHEN 184 => temp2 := 149 ;
		WHEN 185 => temp2 := 55 ;
		WHEN 186 => temp2 := 110 ;
		WHEN 187 => temp2 := 220 ;
		WHEN 188 => temp2 := 165 ;
		WHEN 189 => temp2 := 87 ;
		WHEN 190 => temp2 := 174 ;
		WHEN 191 => temp2 := 65 ;
		WHEN 192 => temp2 := 130 ;
		WHEN 193 => temp2 := 25 ;
		WHEN 194 => temp2 := 50 ;
		WHEN 195 => temp2 := 100 ;
		WHEN 196 => temp2 := 200 ;
		WHEN 197 => temp2 := 141 ;
		WHEN 198 => temp2 := 7 ;
		WHEN 199 => temp2 := 14 ;
		WHEN 200 => temp2 := 28 ;
		WHEN 201 => temp2 := 56 ;
		WHEN 202 => temp2 := 112 ;
		WHEN 203 => temp2 := 224 ;
		WHEN 204 => temp2 := 221 ;
		WHEN 205 => temp2 := 167 ;
		WHEN 206 => temp2 := 83 ;
		WHEN 207 => temp2 := 166 ;
		WHEN 208 => temp2 := 81 ;
		WHEN 209 => temp2 := 162 ;
		WHEN 210 => temp2 := 89 ;
		WHEN 211 => temp2 := 178 ;
		WHEN 212 => temp2 := 121 ;
		WHEN 213 => temp2 := 242 ;
		WHEN 214 => temp2 := 249 ;
		WHEN 215 => temp2 := 239 ;
		WHEN 216 => temp2 := 195 ;
		WHEN 217 => temp2 := 155 ;
		WHEN 218 => temp2 := 43 ;
		WHEN 219 => temp2 := 86 ;
		WHEN 220 => temp2 := 172 ;
		WHEN 221 => temp2 := 69 ;
		WHEN 222 => temp2 := 138 ;
		WHEN 223 => temp2 := 9 ;
		WHEN 224 => temp2 := 18 ;
		WHEN 225 => temp2 := 36 ;
		WHEN 226 => temp2 := 72 ;
		WHEN 227 => temp2 := 144 ;
		WHEN 228 => temp2 := 61 ;
		WHEN 229 => temp2 := 122 ;
		WHEN 230 => temp2 := 244 ;
		WHEN 231 => temp2 := 245 ;
		WHEN 232 => temp2 := 247 ;
		WHEN 233 => temp2 := 243 ;
		WHEN 234 => temp2 := 251 ;
		WHEN 235 => temp2 := 235 ;
		WHEN 236 => temp2 := 203 ;
		WHEN 237 => temp2 := 139 ;
		WHEN 238 => temp2 := 11 ;
		WHEN 239 => temp2 := 22 ;
		WHEN 240 => temp2 := 44 ;
		WHEN 241 => temp2 := 88 ;
		WHEN 242 => temp2 := 176 ;
		WHEN 243 => temp2 := 125 ;
		WHEN 244 => temp2 := 250 ;
		WHEN 245 => temp2 := 233 ;
		WHEN 246 => temp2 := 207 ;
		WHEN 247 => temp2 := 131 ;
		WHEN 248 => temp2 := 27 ;
		WHEN 249 => temp2 := 54 ;
		WHEN 250 => temp2 := 108 ;
		WHEN 251 => temp2 := 216 ;
		WHEN 252 => temp2 := 173 ;
		WHEN 253 => temp2 := 71 ;
		WHEN 254 => temp2 := 142 ;
		WHEN 255 => temp2 := 1 ;
			
		return temp2;
		
		END CASE;
END FUNCTION Convert_to_integer;

end package body my_package;

